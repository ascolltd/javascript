test
podj[pkjvsog
ish;hhd]